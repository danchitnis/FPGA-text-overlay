`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    01:46:38 04/05/2007 
// Design Name: 
// Module Name:    dout_ROM 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module char_ROM(clk, addr, dout);
    input clk;
    input [7:0] addr;
    output [63:0] dout;
	 
	 reg [63:0] dout;
	
	always @(posedge clk)
		case(addr)
			
			
			8'h4A	: // /
						begin
						dout[63:56] 	<= 8'b00000000 ;
						dout[55:48] 	<= 8'b00000011 ;
						dout[47:40] 	<= 8'b00000110 ;
						dout[39:32] 	<=	8'b00001100 ;
						dout[31:24] 	<=	8'b00011000 ;
						dout[23:16]		<=	8'b00110000 ;
						dout[15:8] 		<=	8'b01100000 ;
						dout[7:0]		<=	8'b00000000 ;
						end			
			
			8'h00 : //
						begin
						dout[63:56] 	<= 8'b00000000 ;
						dout[55:48] 	<= 8'b00000000 ;
						dout[47:40] 	<= 8'b00000000 ;
						dout[39:32] 	<=	8'b00000000 ;
						dout[31:24] 	<=	8'b00000000 ;
						dout[23:16]		<=	8'b00000000 ;
						dout[15:8] 		<=	8'b00000000 ;
						dout[7:0]		<=	8'b00000000 ;
						end
						
	
						
			8'h16	: 	//1
						begin
						dout[63:56]		<= 8'b00011000 ;
						dout[55:48]		<= 8'b00011000 ;
						dout[47:40]		<= 8'b00111000 ;
						dout[39:32]		<=	8'b00011000 ;
						dout[31:24]		<=	8'b00011000 ;
						dout[23:16]		<=	8'b00011000 ;
						dout[15:8]		<=	8'b01111110 ;
						dout[7:0]		<=	8'b00000000 ;
						end
						
			8'hFF	:	//
						begin
						dout[63:56] 	<= 8'b01111110 ;
						dout[55:48] 	<= 8'b01111110 ;
						dout[47:40] 	<= 8'b01111110 ;
						dout[39:32] 	<=	8'b01111110 ;
						dout[31:24] 	<=	8'b01111110 ;
						dout[23:16]		<=	8'b01111110 ;
						dout[15:8] 		<=	8'b01111110 ;
						dout[7:0]		<=	8'b00000000 ;
						end
						
							
			8'h1E	:	//2
						begin
						dout[63:56]		<= 8'b00111100 ;
						dout[55:48]		<= 8'b01100110 ;
						dout[47:40]		<= 8'b00000110 ;
						dout[39:32]		<=	8'b00001100 ;
						dout[31:24]		<=	8'b00110000 ;
						dout[23:16]		<=	8'b01100000 ;
						dout[15:8] 		<=	8'b01111110 ;
						dout[7:0]		<=	8'b00000000 ;
						end
						
												
			8'h26	:	//3
						begin
						dout[63:56]		<= 8'b00111100 ;
						dout[55:48] 	<= 8'b01100110 ;
						dout[47:40] 	<= 8'b00000110 ;
						dout[39:32]		<=	8'b00011100 ;
						dout[31:24] 	<=	8'b00000110 ;
						dout[23:16]		<=	8'b01100110 ;
						dout[15:8] 		<=	8'b00111100 ;
						dout[7:0]		<=	8'b00000000 ;
						end
						
			8'h25	: //4
						begin
						dout[63:56]		<= 8'b00000110 ;
						dout[55:48]		<= 8'b00001110 ;
						dout[47:40]		<= 8'b00011110 ;
						dout[39:32] 	<=	8'b01100110 ;
						dout[31:24] 	<=	8'b01111111 ;
						dout[23:16]		<=	8'b00000110 ;
						dout[15:8]		<=	8'b00000110 ;
						dout[7:0]		<=	8'b00000000 ;
						end
	 
			8'h2E	: // 5
						begin
						dout[63:56] 	<= 8'b01111110 ;
						dout[55:48] 	<= 8'b01100000 ;
						dout[47:40] 	<= 8'b01111100 ;
						dout[39:32] 	<=	8'b00000110 ;
						dout[31:24] 	<=	8'b00000110 ;
						dout[23:16]		<=	8'b01100110 ;
						dout[15:8] 		<=	8'b00111100 ;
						dout[7:0]		<=	8'b00000000 ;
						end


			8'h36	: // 6
						begin
						dout[63:56] 	<= 8'b00111100 ;
						dout[55:48] 	<= 8'b01100110 ;
						dout[47:40] 	<= 8'b01100000 ;
						dout[39:32] 	<=	8'b01111100 ;
						dout[31:24] 	<=	8'b01100110 ;
						dout[23:16]		<=	8'b01100110 ;
						dout[15:8] 		<=	8'b00111100 ;
						dout[7:0]		<=	8'b00000000 ;
						end
						

			8'h3D	: // 7
						begin
						dout[63:56] 	<= 8'b01111110 ;
						dout[55:48] 	<= 8'b01100110 ;
						dout[47:40] 	<= 8'b00001100 ;
						dout[39:32] 	<=	8'b00011000 ;
						dout[31:24] 	<=	8'b00011000 ;
						dout[23:16]		<=	8'b00011000 ;
						dout[15:8] 		<=	8'b00011000 ;
						dout[7:0]		<=	8'b00000000 ;
						end	
				
			8'h3E	: // 8
						begin
						dout[63:56] 	<= 8'b00111100 ;
						dout[55:48] 	<= 8'b01100110 ;
						dout[47:40] 	<= 8'b01100110 ;
						dout[39:32] 	<=	8'b00111100 ;
						dout[31:24] 	<=	8'b01100110 ;
						dout[23:16]		<=	8'b01100110 ;
						dout[15:8] 		<=	8'b00111100 ;
						dout[7:0]		<=	8'b00000000 ;
						end
 
			8'h46	: // 9
						begin
						dout[63:56] 	<= 8'b00111100 ;
						dout[55:48] 	<= 8'b01100110 ;
						dout[47:40] 	<= 8'b01100110 ;
						dout[39:32] 	<=	8'b00111110 ;
						dout[31:24] 	<=	8'b00000110 ;
						dout[23:16]		<=	8'b01100110 ;
						dout[15:8] 		<=	8'b00111100 ;
						dout[7:0]		<=	8'b00000000 ;
						end
			8'h49	: // .
						begin
						dout[63:56] 	<= 8'b00000000 ;
						dout[55:48] 	<= 8'b00000000 ;
						dout[47:40] 	<= 8'b00000000 ;
						dout[39:32] 	<=	8'b00000000 ;
						dout[31:24] 	<=	8'b00000000 ;
						dout[23:16]		<=	8'b00011000 ;
						dout[15:8] 		<=	8'b00011000 ;
						dout[7:0]		<=	8'b00000000 ;
						end

			
	
			8'h45	: // 0
						begin
						dout[63:56] 	<= 8'b00111100 ;
						dout[55:48] 	<= 8'b01100110 ;
						dout[47:40] 	<= 8'b01101110 ;
						dout[39:32] 	<=	8'b01110110 ;
						dout[31:24] 	<=	8'b01100110 ;
						dout[23:16]		<=	8'b01100110 ;
						dout[15:8] 		<=	8'b00111100 ;
						dout[7:0]		<=	8'b00000000 ;
						end
						
			/*8'h	: // :
						begin
						dout[63:56] 	<= 8'b00000000 ;
						dout[55:48] 	<= 8'b00011000 ;
						dout[47:40] 	<= 8'b00011000 ;
						dout[39:32] 	<=	8'b00000000 ;
						dout[31:24] 	<=	8'b00011000 ;
						dout[23:16]		<=	8'b00011000 ;
						dout[15:8] 		<=	8'b00000000 ;
						dout[7:0]		<=	8'b00000000 ;
						end*/
						
			8'h4C	: // ;
						begin
						dout[63:56] 	<= 8'b00000000 ;
						dout[55:48] 	<= 8'b00011000 ;
						dout[47:40] 	<= 8'b00011000 ;
						dout[39:32] 	<=	8'b00000000 ;
						dout[31:24] 	<=	8'b00011000 ;
						dout[23:16]		<=	8'b00011000 ;
						dout[15:8] 		<=	8'b00110000 ;
						dout[7:0]		<=	8'b00000000 ;
						end
						
			8'h1C	: //A
						begin
						dout[63:56] 	<= 8'b00011000 ;
						dout[55:48] 	<= 8'b00111100 ;
						dout[47:40] 	<= 8'b01100110 ;
						dout[39:32] 	<=	8'b01111110 ;
						dout[31:24] 	<=	8'b01100110 ;
						dout[23:16]		<=	8'b01100110 ;
						dout[15:8] 		<=	8'b01100110 ;
						dout[7:0]		<=	8'b00000000 ;
						end

			8'h32	: // B
						begin
						dout[63:56] 	<= 8'b01111100 ;
						dout[55:48] 	<= 8'b01100110 ;
						dout[47:40] 	<= 8'b01100110 ;
						dout[39:32] 	<=	8'b01111100 ;
						dout[31:24] 	<=	8'b01100110 ;
						dout[23:16]		<=	8'b01100110 ;
						dout[15:8] 		<=	8'b01111100 ;
						dout[7:0]		<=	8'b00000000 ;
						end
						
			8'h21	: // C
						begin
						dout[63:56] 	<= 8'b00111100 ;
						dout[55:48] 	<= 8'b01100110 ;
						dout[47:40] 	<= 8'b01100000 ;
						dout[39:32] 	<=	8'b01100000 ;
						dout[31:24] 	<=	8'b01100000 ;
						dout[23:16]		<=	8'b01100110 ;
						dout[15:8] 		<=	8'b00111100 ;
						dout[7:0]		<=	8'b00000000 ;
						end
						
			8'h23	: // D
						begin
						dout[63:56] 	<= 8'b01111000 ;
						dout[55:48] 	<= 8'b01101100 ;
						dout[47:40] 	<= 8'b01100110 ;
						dout[39:32] 	<=	8'b01100110 ;
						dout[31:24] 	<=	8'b01100110 ;
						dout[23:16]		<=	8'b01101100 ;
						dout[15:8] 		<=	8'b01111000 ;
						dout[7:0]		<=	8'b00000000 ;
						end
						
			8'h24	: // E
						begin
						dout[63:56] 	<= 8'b01111110 ;
						dout[55:48] 	<= 8'b01100000 ;
						dout[47:40] 	<= 8'b01100000 ;
						dout[39:32] 	<=	8'b01111000 ;
						dout[31:24] 	<=	8'b01100000 ;
						dout[23:16]		<=	8'b01100000 ;
						dout[15:8] 		<=	8'b01111110 ;
						dout[7:0]		<=	8'b00000000 ;
						end
						
			8'h2B	: // F
						begin
						dout[63:56] 	<= 8'b01111110 ;
						dout[55:48] 	<= 8'b01100000 ;
						dout[47:40] 	<= 8'b01100000 ;
						dout[39:32] 	<=	8'b01111000 ;
						dout[31:24] 	<=	8'b01100000 ;
						dout[23:16]		<=	8'b01100000 ;
						dout[15:8] 		<=	8'b01100000 ;
						dout[7:0]		<=	8'b00000000 ;
						end
						
			8'h34	: // G
						begin
						dout[63:56] 	<= 8'b00111100 ;
						dout[55:48] 	<= 8'b01100110 ;
						dout[47:40] 	<= 8'b01100000 ;
						dout[39:32] 	<=	8'b01101110 ;
						dout[31:24] 	<=	8'b01100110 ;
						dout[23:16]		<=	8'b01100110 ;
						dout[15:8] 		<=	8'b00111100 ;
						dout[7:0]		<=	8'b00000000 ;
						end
						
			8'h33	: // H
						begin
						dout[63:56] 	<= 8'b01100110 ;
						dout[55:48] 	<= 8'b01100110 ;
						dout[47:40] 	<= 8'b01100110 ;
						dout[39:32] 	<=	8'b01111110 ;
						dout[31:24] 	<=	8'b01100110 ;
						dout[23:16]		<=	8'b01100110 ;
						dout[15:8] 		<=	8'b01100110 ;
						dout[7:0]		<=	8'b00000000 ;
						end
						
			8'h43	: // I
						begin
						dout[63:56] 	<= 8'b00111100 ;
						dout[55:48] 	<= 8'b00011000 ;
						dout[47:40] 	<= 8'b00011000 ;
						dout[39:32] 	<=	8'b00011000 ;
						dout[31:24] 	<=	8'b00011000 ;
						dout[23:16]		<=	8'b00011000 ;
						dout[15:8] 		<=	8'b00111100 ;
						dout[7:0]		<=	8'b00000000 ;
						end
						
			8'h3B	: // J
						begin
						dout[63:56] 	<= 8'b00011110 ;
						dout[55:48] 	<= 8'b00001100 ;
						dout[47:40] 	<= 8'b00001100 ;
						dout[39:32] 	<=	8'b00001100 ;
						dout[31:24] 	<=	8'b00001100 ;
						dout[23:16]		<=	8'b01101100 ;
						dout[15:8] 		<=	8'b00111000 ;
						dout[7:0]		<=	8'b00000000 ;
						end
						
			8'h42	: // K
						begin
						dout[63:56] 	<= 8'b01100110 ;
						dout[55:48] 	<= 8'b01101100 ;
						dout[47:40] 	<= 8'b01111000 ;
						dout[39:32] 	<=	8'b01110000 ;
						dout[31:24] 	<=	8'b01111000 ;
						dout[23:16]		<=	8'b01101100 ;
						dout[15:8] 		<=	8'b01100110 ;
						dout[7:0]		<=	8'b00000000 ;
						end
						
			8'h4B	: // L
						begin
						dout[63:56] 	<= 8'b01100000 ;
						dout[55:48] 	<= 8'b01100000 ;
						dout[47:40] 	<= 8'b01100000 ;
						dout[39:32] 	<=	8'b01100000 ;
						dout[31:24] 	<=	8'b01100000 ;
						dout[23:16]		<=	8'b01100000 ;
						dout[15:8] 		<=	8'b01111110 ;
						dout[7:0]		<=	8'b00000000 ;
						end
						
			8'h3A	: // M
						begin
						dout[63:56] 	<= 8'b01100011 ;
						dout[55:48] 	<= 8'b01110111 ;
						dout[47:40] 	<= 8'b01111111 ;
						dout[39:32] 	<=	8'b01101011 ;
						dout[31:24] 	<=	8'b01100011 ;
						dout[23:16]		<=	8'b01100011 ;
						dout[15:8] 		<=	8'b01100011 ;
						dout[7:0]		<=	8'b00000000 ;
						end
						
			8'h31	: // N
						begin
						dout[63:56] 	<= 8'b01100110 ;
						dout[55:48] 	<= 8'b01110110 ;
						dout[47:40] 	<= 8'b01111110 ;
						dout[39:32] 	<=	8'b01111110 ;
						dout[31:24] 	<=	8'b01101110 ;
						dout[23:16]		<=	8'b01100110 ;
						dout[15:8] 		<=	8'b01100110 ;
						dout[7:0]		<=	8'b00000000 ;
						end
						
			8'h44	: // O
						begin
						dout[63:56] 	<= 8'b00111100 ;
						dout[55:48] 	<= 8'b01100110 ;
						dout[47:40] 	<= 8'b01100110 ;
						dout[39:32] 	<=	8'b01100110 ;
						dout[31:24] 	<=	8'b01100110 ;
						dout[23:16]		<=	8'b01100110 ;
						dout[15:8] 		<=	8'b00111100 ;
						dout[7:0]		<=	8'b00000000 ;
						end
						
			8'h4D	: // P
						begin
						dout[63:56] 	<= 8'b01111100 ;
						dout[55:48] 	<= 8'b01100110 ;
						dout[47:40] 	<= 8'b01100110 ;
						dout[39:32] 	<=	8'b01111100 ;
						dout[31:24] 	<=	8'b01100000 ;
						dout[23:16]		<=	8'b01100000 ;
						dout[15:8] 		<=	8'b01100000 ;
						dout[7:0]		<=	8'b00000000 ;
						end
						
			8'h15	: // Q
						begin
						dout[63:56] 	<= 8'b00111100 ;
						dout[55:48] 	<= 8'b01100110 ;
						dout[47:40] 	<= 8'b01100110 ;
						dout[39:32] 	<=	8'b01100110 ;
						dout[31:24] 	<=	8'b01100110 ;
						dout[23:16]		<=	8'b00111100 ;
						dout[15:8] 		<=	8'b00001110 ;
						dout[7:0]		<=	8'b00000000 ;
						end
						
			8'h2D	: // R
						begin
						dout[63:56] 	<= 8'b01111100 ;
						dout[55:48] 	<= 8'b01100110 ;
						dout[47:40] 	<= 8'b01100110 ;
						dout[39:32] 	<=	8'b01111100 ;
						dout[31:24] 	<=	8'b01111000 ;
						dout[23:16]		<=	8'b01101100 ;
						dout[15:8] 		<=	8'b01100110 ;
						dout[7:0]		<=	8'b00000000 ;
						end
						
			8'h1B	: // S
						begin
						dout[63:56] 	<= 8'b00111100 ;
						dout[55:48] 	<= 8'b01100110 ;
						dout[47:40] 	<= 8'b01100000 ;
						dout[39:32] 	<=	8'b00111100 ;
						dout[31:24] 	<=	8'b00000110 ;
						dout[23:16]		<=	8'b01100110 ;
						dout[15:8] 		<=	8'b00111100 ;
						dout[7:0]		<=	8'b00000000 ;
						end
						
			8'h2C	: //T
						begin
						dout[63:56] 	<= 8'b01111110 ;
						dout[55:48] 	<= 8'b00011000 ;
						dout[47:40] 	<= 8'b00011000 ;
						dout[39:32] 	<=	8'b00011000 ;
						dout[31:24] 	<=	8'b00011000 ;
						dout[23:16]		<=	8'b00011000 ;
						dout[15:8] 		<=	8'b00011000 ;
						dout[7:0]		<=	8'b00000000 ;
						end
						
			8'h3C	: //U
						begin
						dout[63:56] 	<= 8'b01100110 ;
						dout[55:48] 	<= 8'b01100110 ;
						dout[47:40] 	<= 8'b01100110 ;
						dout[39:32] 	<=	8'b01100110 ;
						dout[31:24] 	<=	8'b01100110 ;
						dout[23:16]		<=	8'b01100110 ;
						dout[15:8] 		<=	8'b00111100 ;
						dout[7:0]		<=	8'b00000000 ;
						end
						
			8'h2A	: //V
						begin
						dout[63:56] 	<= 8'b01100110 ;
						dout[55:48] 	<= 8'b01100110 ;
						dout[47:40] 	<= 8'b01100110 ;
						dout[39:32] 	<=	8'b01100110 ;
						dout[31:24] 	<=	8'b01100110 ;
						dout[23:16]		<=	8'b00111100 ;
						dout[15:8] 		<=	8'b00011000 ;
						dout[7:0]		<=	8'b00000000 ;
						end
						
			8'h1D	: //W
						begin
						dout[63:56] 	<= 8'b01100011 ;
						dout[55:48] 	<= 8'b01100011 ;
						dout[47:40] 	<= 8'b01100011 ;
						dout[39:32] 	<=	8'b01101011 ;
						dout[31:24] 	<=	8'b01111111 ;
						dout[23:16]		<=	8'b01110111 ;
						dout[15:8] 		<=	8'b01100011 ;
						dout[7:0]		<=	8'b00000000 ;
						end
						
			8'h22	: //X
						begin
						dout[63:56] 	<= 8'b01100110 ;
						dout[55:48] 	<= 8'b01100110 ;
						dout[47:40] 	<= 8'b00111100 ;
						dout[39:32] 	<=	8'b00011000 ;
						dout[31:24] 	<=	8'b00111100 ;
						dout[23:16]		<=	8'b01100110 ;
						dout[15:8] 		<=	8'b01100110 ;
						dout[7:0]		<=	8'b00000000 ;
						end
						
			8'h35	: //Y
						begin
						dout[63:56] 	<= 8'b01100110 ;
						dout[55:48] 	<= 8'b01100110 ;
						dout[47:40] 	<= 8'b01100110 ;
						dout[39:32] 	<=	8'b00111100 ;
						dout[31:24] 	<=	8'b00011000 ;
						dout[23:16]		<=	8'b00011000 ;
						dout[15:8] 		<=	8'b00011000 ;
						dout[7:0]		<=	8'b00000000 ;
						end
						
			/*8'h	: //
						begin
						dout[63:56] 	<= 8'b ;
						dout[55:48] 	<= 8'b ;
						dout[47:40] 	<= 8'b ;
						dout[39:32] 	<=	8'b ;
						dout[31:24] 	<=	8'b ;
						dout[23:16]		<=	8'b ;
						dout[15:8] 		<=	8'b ;
						dout[7:0]		<=	8'b00000000 ;
						end*/
						
			8'h1A	: // Z
						begin
						dout[63:56] 	<= 8'b01111110 ;
						dout[55:48] 	<= 8'b00000110 ;
						dout[47:40] 	<= 8'b00001100 ;
						dout[39:32] 	<=	8'b00011000 ;
						dout[31:24] 	<=	8'b00110000 ;
						dout[23:16]		<=	8'b01100000 ;
						dout[15:8] 		<=	8'b01111110 ;
						dout[7:0]		<=	8'b00000000 ;
						end
			
			default dout<=0;
			
		endcase

endmodule
